module LolaP_round_w
(
    input [256:0] round_i,
    output [256:0] round_o
);

wire [256:0] after_pi_s;
wire [256:0] after_theta_s;

// Pi step
generate
    genvar gen_j;
    for (gen_j = 0; gen_j < 257; gen_j = gen_j + 1) begin: pi_step
        assign after_pi_s[gen_j] = round_i[(121*gen_j) % 257];
    end
endgenerate

// Theta and iota steps
assign after_theta_s[12]  = after_pi_s[12]  ^ after_pi_s[15]  ^ after_pi_s[22];  
assign after_theta_s[56]  = after_pi_s[56]  ^ after_pi_s[59]  ^ after_pi_s[66]; 
assign after_theta_s[90]  = after_pi_s[90]  ^ after_pi_s[93]  ^ after_pi_s[100];
assign after_theta_s[163] = after_pi_s[163] ^ after_pi_s[166] ^ after_pi_s[173];
assign after_theta_s[161] = after_pi_s[161] ^ after_pi_s[164] ^ after_pi_s[171];
assign after_theta_s[66]  = after_pi_s[66]  ^ after_pi_s[69]  ^ after_pi_s[76];
assign after_theta_s[51]  = after_pi_s[51]  ^ after_pi_s[54]  ^ after_pi_s[61];
assign after_theta_s[238] = after_pi_s[238] ^ after_pi_s[241] ^ after_pi_s[248];
assign after_theta_s[254] = after_pi_s[254] ^ after_pi_s[0]   ^ after_pi_s[7];
assign after_theta_s[243] = after_pi_s[243] ^ after_pi_s[246] ^ after_pi_s[253];
assign after_theta_s[106] = after_pi_s[106] ^ after_pi_s[109] ^ after_pi_s[116];
assign after_theta_s[152] = after_pi_s[152] ^ after_pi_s[155] ^ after_pi_s[162];
assign after_theta_s[24]  = after_pi_s[24]  ^ after_pi_s[27]  ^ after_pi_s[34];
assign after_theta_s[112] = after_pi_s[112] ^ after_pi_s[115] ^ after_pi_s[122];
assign after_theta_s[180] = after_pi_s[180] ^ after_pi_s[183] ^ after_pi_s[190];
assign after_theta_s[69]  = after_pi_s[69]  ^ after_pi_s[72]  ^ after_pi_s[79];
assign after_theta_s[65]  = after_pi_s[65]  ^ after_pi_s[68]  ^ after_pi_s[75];
assign after_theta_s[132] = after_pi_s[132] ^ after_pi_s[135] ^ after_pi_s[142];
assign after_theta_s[102] = after_pi_s[102] ^ after_pi_s[105] ^ after_pi_s[112];
assign after_theta_s[219] = after_pi_s[219] ^ after_pi_s[222] ^ after_pi_s[229];
assign after_theta_s[251] = after_pi_s[251] ^ after_pi_s[254] ^ after_pi_s[4];
assign after_theta_s[229] = after_pi_s[229] ^ after_pi_s[232] ^ after_pi_s[239];
assign after_theta_s[212] = after_pi_s[212] ^ after_pi_s[215] ^ after_pi_s[222];
assign after_theta_s[47]  = after_pi_s[47]  ^ after_pi_s[50]  ^ after_pi_s[57];
assign after_theta_s[48]  = after_pi_s[48]  ^ after_pi_s[51]  ^ after_pi_s[58];
assign after_theta_s[224] = after_pi_s[224] ^ after_pi_s[227] ^ after_pi_s[234];
assign after_theta_s[103] = after_pi_s[103] ^ after_pi_s[106] ^ after_pi_s[113];
assign after_theta_s[138] = after_pi_s[138] ^ after_pi_s[141] ^ after_pi_s[148];
assign after_theta_s[130] = after_pi_s[130] ^ after_pi_s[133] ^ after_pi_s[140];
assign after_theta_s[7]   = after_pi_s[7]   ^ after_pi_s[10]  ^ after_pi_s[17];
assign after_theta_s[204] = after_pi_s[204] ^ after_pi_s[207] ^ after_pi_s[214];
assign after_theta_s[181] = after_pi_s[181] ^ after_pi_s[184] ^ after_pi_s[191];
assign after_theta_s[245] = after_pi_s[245] ^ after_pi_s[248] ^ after_pi_s[255];
assign after_theta_s[0] = ~(after_pi_s[0] ^ after_pi_s[3] ^ after_pi_s[10]);
assign after_theta_s[36] = after_pi_s[36] ^ after_pi_s[39] ^ after_pi_s[46];
assign after_theta_s[60] = after_pi_s[60] ^ after_pi_s[63] ^ after_pi_s[70];
assign after_theta_s[72] = after_pi_s[72] ^ after_pi_s[75] ^ after_pi_s[82];
assign after_theta_s[84] = after_pi_s[84] ^ after_pi_s[87] ^ after_pi_s[94];
assign after_theta_s[96] = after_pi_s[96] ^ after_pi_s[99] ^ after_pi_s[106];
assign after_theta_s[108] = after_pi_s[108] ^ after_pi_s[111] ^ after_pi_s[118];
assign after_theta_s[120] = after_pi_s[120] ^ after_pi_s[123] ^ after_pi_s[130];
assign after_theta_s[144] = after_pi_s[144] ^ after_pi_s[147] ^ after_pi_s[154];
assign after_theta_s[156] = after_pi_s[156] ^ after_pi_s[159] ^ after_pi_s[166];
assign after_theta_s[168] = after_pi_s[168] ^ after_pi_s[171] ^ after_pi_s[178];
assign after_theta_s[192] = after_pi_s[192] ^ after_pi_s[195] ^ after_pi_s[202];
assign after_theta_s[216] = after_pi_s[216] ^ after_pi_s[219] ^ after_pi_s[226];
assign after_theta_s[228] = after_pi_s[228] ^ after_pi_s[231] ^ after_pi_s[238];
assign after_theta_s[240] = after_pi_s[240] ^ after_pi_s[243] ^ after_pi_s[250];
assign after_theta_s[252] = after_pi_s[252] ^ after_pi_s[255] ^ after_pi_s[5];
assign after_theta_s[19] = after_pi_s[19] ^ after_pi_s[22] ^ after_pi_s[29];
assign after_theta_s[31] = after_pi_s[31] ^ after_pi_s[34] ^ after_pi_s[41];
assign after_theta_s[43] = after_pi_s[43] ^ after_pi_s[46] ^ after_pi_s[53];
assign after_theta_s[55] = after_pi_s[55] ^ after_pi_s[58] ^ after_pi_s[65];
assign after_theta_s[67] = after_pi_s[67] ^ after_pi_s[70] ^ after_pi_s[77];
assign after_theta_s[79] = after_pi_s[79] ^ after_pi_s[82] ^ after_pi_s[89];
assign after_theta_s[91] = after_pi_s[91] ^ after_pi_s[94] ^ after_pi_s[101];
assign after_theta_s[115] = after_pi_s[115] ^ after_pi_s[118] ^ after_pi_s[125];
assign after_theta_s[127] = after_pi_s[127] ^ after_pi_s[130] ^ after_pi_s[137];
assign after_theta_s[139] = after_pi_s[139] ^ after_pi_s[142] ^ after_pi_s[149];
assign after_theta_s[151] = after_pi_s[151] ^ after_pi_s[154] ^ after_pi_s[161];
assign after_theta_s[175] = after_pi_s[175] ^ after_pi_s[178] ^ after_pi_s[185];
assign after_theta_s[187] = after_pi_s[187] ^ after_pi_s[190] ^ after_pi_s[197];
assign after_theta_s[199] = after_pi_s[199] ^ after_pi_s[202] ^ after_pi_s[209];
assign after_theta_s[211] = after_pi_s[211] ^ after_pi_s[214] ^ after_pi_s[221];
assign after_theta_s[223] = after_pi_s[223] ^ after_pi_s[226] ^ after_pi_s[233];
assign after_theta_s[235] = after_pi_s[235] ^ after_pi_s[238] ^ after_pi_s[245];
assign after_theta_s[247] = after_pi_s[247] ^ after_pi_s[250] ^ after_pi_s[0];
assign after_theta_s[2] = after_pi_s[2] ^ after_pi_s[5] ^ after_pi_s[12];
assign after_theta_s[14] = after_pi_s[14] ^ after_pi_s[17] ^ after_pi_s[24];
assign after_theta_s[26] = after_pi_s[26] ^ after_pi_s[29] ^ after_pi_s[36];
assign after_theta_s[38] = after_pi_s[38] ^ after_pi_s[41] ^ after_pi_s[48];
assign after_theta_s[50] = after_pi_s[50] ^ after_pi_s[53] ^ after_pi_s[60];
assign after_theta_s[62] = after_pi_s[62] ^ after_pi_s[65] ^ after_pi_s[72];
assign after_theta_s[74] = after_pi_s[74] ^ after_pi_s[77] ^ after_pi_s[84];
assign after_theta_s[86] = after_pi_s[86] ^ after_pi_s[89] ^ after_pi_s[96];
assign after_theta_s[98] = after_pi_s[98] ^ after_pi_s[101] ^ after_pi_s[108];
assign after_theta_s[110] = after_pi_s[110] ^ after_pi_s[113] ^ after_pi_s[120];
assign after_theta_s[122] = after_pi_s[122] ^ after_pi_s[125] ^ after_pi_s[132];
assign after_theta_s[134] = after_pi_s[134] ^ after_pi_s[137] ^ after_pi_s[144];
assign after_theta_s[146] = after_pi_s[146] ^ after_pi_s[149] ^ after_pi_s[156];
assign after_theta_s[158] = after_pi_s[158] ^ after_pi_s[161] ^ after_pi_s[168];
assign after_theta_s[170] = after_pi_s[170] ^ after_pi_s[173] ^ after_pi_s[180];
assign after_theta_s[182] = after_pi_s[182] ^ after_pi_s[185] ^ after_pi_s[192];
assign after_theta_s[194] = after_pi_s[194] ^ after_pi_s[197] ^ after_pi_s[204];
assign after_theta_s[206] = after_pi_s[206] ^ after_pi_s[209] ^ after_pi_s[216];
assign after_theta_s[218] = after_pi_s[218] ^ after_pi_s[221] ^ after_pi_s[228];
assign after_theta_s[230] = after_pi_s[230] ^ after_pi_s[233] ^ after_pi_s[240];
assign after_theta_s[242] = after_pi_s[242] ^ after_pi_s[245] ^ after_pi_s[252];
assign after_theta_s[9] = after_pi_s[9] ^ after_pi_s[12] ^ after_pi_s[19];
assign after_theta_s[21] = after_pi_s[21] ^ after_pi_s[24] ^ after_pi_s[31];
assign after_theta_s[33] = after_pi_s[33] ^ after_pi_s[36] ^ after_pi_s[43];
assign after_theta_s[45] = after_pi_s[45] ^ after_pi_s[48] ^ after_pi_s[55];
assign after_theta_s[57] = after_pi_s[57] ^ after_pi_s[60] ^ after_pi_s[67];
assign after_theta_s[81] = after_pi_s[81] ^ after_pi_s[84] ^ after_pi_s[91];
assign after_theta_s[93] = after_pi_s[93] ^ after_pi_s[96] ^ after_pi_s[103];
assign after_theta_s[105] = after_pi_s[105] ^ after_pi_s[108] ^ after_pi_s[115];
assign after_theta_s[117] = after_pi_s[117] ^ after_pi_s[120] ^ after_pi_s[127];
assign after_theta_s[129] = after_pi_s[129] ^ after_pi_s[132] ^ after_pi_s[139];
assign after_theta_s[141] = after_pi_s[141] ^ after_pi_s[144] ^ after_pi_s[151];
assign after_theta_s[153] = after_pi_s[153] ^ after_pi_s[156] ^ after_pi_s[163];
assign after_theta_s[165] = after_pi_s[165] ^ after_pi_s[168] ^ after_pi_s[175];
assign after_theta_s[177] = after_pi_s[177] ^ after_pi_s[180] ^ after_pi_s[187];
assign after_theta_s[189] = after_pi_s[189] ^ after_pi_s[192] ^ after_pi_s[199];
assign after_theta_s[201] = after_pi_s[201] ^ after_pi_s[204] ^ after_pi_s[211];
assign after_theta_s[213] = after_pi_s[213] ^ after_pi_s[216] ^ after_pi_s[223];
assign after_theta_s[225] = after_pi_s[225] ^ after_pi_s[228] ^ after_pi_s[235];
assign after_theta_s[237] = after_pi_s[237] ^ after_pi_s[240] ^ after_pi_s[247];
assign after_theta_s[249] = after_pi_s[249] ^ after_pi_s[252] ^ after_pi_s[2];
assign after_theta_s[4] = after_pi_s[4] ^ after_pi_s[7] ^ after_pi_s[14];
assign after_theta_s[16] = after_pi_s[16] ^ after_pi_s[19] ^ after_pi_s[26];
assign after_theta_s[28] = after_pi_s[28] ^ after_pi_s[31] ^ after_pi_s[38];
assign after_theta_s[40] = after_pi_s[40] ^ after_pi_s[43] ^ after_pi_s[50];
assign after_theta_s[52] = after_pi_s[52] ^ after_pi_s[55] ^ after_pi_s[62];
assign after_theta_s[64] = after_pi_s[64] ^ after_pi_s[67] ^ after_pi_s[74];
assign after_theta_s[76] = after_pi_s[76] ^ after_pi_s[79] ^ after_pi_s[86];
assign after_theta_s[88] = after_pi_s[88] ^ after_pi_s[91] ^ after_pi_s[98];
assign after_theta_s[100] = after_pi_s[100] ^ after_pi_s[103] ^ after_pi_s[110];
assign after_theta_s[124] = after_pi_s[124] ^ after_pi_s[127] ^ after_pi_s[134];
assign after_theta_s[136] = after_pi_s[136] ^ after_pi_s[139] ^ after_pi_s[146];
assign after_theta_s[148] = after_pi_s[148] ^ after_pi_s[151] ^ after_pi_s[158];
assign after_theta_s[160] = after_pi_s[160] ^ after_pi_s[163] ^ after_pi_s[170];
assign after_theta_s[172] = after_pi_s[172] ^ after_pi_s[175] ^ after_pi_s[182];
assign after_theta_s[184] = after_pi_s[184] ^ after_pi_s[187] ^ after_pi_s[194];
assign after_theta_s[196] = after_pi_s[196] ^ after_pi_s[199] ^ after_pi_s[206];
assign after_theta_s[208] = after_pi_s[208] ^ after_pi_s[211] ^ after_pi_s[218];
assign after_theta_s[220] = after_pi_s[220] ^ after_pi_s[223] ^ after_pi_s[230];
assign after_theta_s[232] = after_pi_s[232] ^ after_pi_s[235] ^ after_pi_s[242];
assign after_theta_s[244] = after_pi_s[244] ^ after_pi_s[247] ^ after_pi_s[254];
assign after_theta_s[256] = after_pi_s[256] ^ after_pi_s[2] ^ after_pi_s[9];
assign after_theta_s[11] = after_pi_s[11] ^ after_pi_s[14] ^ after_pi_s[21];
assign after_theta_s[23] = after_pi_s[23] ^ after_pi_s[26] ^ after_pi_s[33];
assign after_theta_s[35] = after_pi_s[35] ^ after_pi_s[38] ^ after_pi_s[45];
assign after_theta_s[59] = after_pi_s[59] ^ after_pi_s[62] ^ after_pi_s[69];
assign after_theta_s[71] = after_pi_s[71] ^ after_pi_s[74] ^ after_pi_s[81];
assign after_theta_s[83] = after_pi_s[83] ^ after_pi_s[86] ^ after_pi_s[93];
assign after_theta_s[95] = after_pi_s[95] ^ after_pi_s[98] ^ after_pi_s[105];
assign after_theta_s[107] = after_pi_s[107] ^ after_pi_s[110] ^ after_pi_s[117];
assign after_theta_s[119] = after_pi_s[119] ^ after_pi_s[122] ^ after_pi_s[129];
assign after_theta_s[131] = after_pi_s[131] ^ after_pi_s[134] ^ after_pi_s[141];
assign after_theta_s[143] = after_pi_s[143] ^ after_pi_s[146] ^ after_pi_s[153];
assign after_theta_s[155] = after_pi_s[155] ^ after_pi_s[158] ^ after_pi_s[165];
assign after_theta_s[167] = after_pi_s[167] ^ after_pi_s[170] ^ after_pi_s[177];
assign after_theta_s[179] = after_pi_s[179] ^ after_pi_s[182] ^ after_pi_s[189];
assign after_theta_s[191] = after_pi_s[191] ^ after_pi_s[194] ^ after_pi_s[201];
assign after_theta_s[203] = after_pi_s[203] ^ after_pi_s[206] ^ after_pi_s[213];
assign after_theta_s[215] = after_pi_s[215] ^ after_pi_s[218] ^ after_pi_s[225];
assign after_theta_s[227] = after_pi_s[227] ^ after_pi_s[230] ^ after_pi_s[237];
assign after_theta_s[239] = after_pi_s[239] ^ after_pi_s[242] ^ after_pi_s[249];
assign after_theta_s[6] = after_pi_s[6] ^ after_pi_s[9] ^ after_pi_s[16];
assign after_theta_s[18] = after_pi_s[18] ^ after_pi_s[21] ^ after_pi_s[28];
assign after_theta_s[30] = after_pi_s[30] ^ after_pi_s[33] ^ after_pi_s[40];
assign after_theta_s[42] = after_pi_s[42] ^ after_pi_s[45] ^ after_pi_s[52];
assign after_theta_s[54] = after_pi_s[54] ^ after_pi_s[57] ^ after_pi_s[64];
assign after_theta_s[78] = after_pi_s[78] ^ after_pi_s[81] ^ after_pi_s[88];
assign after_theta_s[114] = after_pi_s[114] ^ after_pi_s[117] ^ after_pi_s[124];
assign after_theta_s[126] = after_pi_s[126] ^ after_pi_s[129] ^ after_pi_s[136];
assign after_theta_s[150] = after_pi_s[150] ^ after_pi_s[153] ^ after_pi_s[160];
assign after_theta_s[162] = after_pi_s[162] ^ after_pi_s[165] ^ after_pi_s[172];
assign after_theta_s[174] = after_pi_s[174] ^ after_pi_s[177] ^ after_pi_s[184];
assign after_theta_s[186] = after_pi_s[186] ^ after_pi_s[189] ^ after_pi_s[196];
assign after_theta_s[198] = after_pi_s[198] ^ after_pi_s[201] ^ after_pi_s[208];
assign after_theta_s[210] = after_pi_s[210] ^ after_pi_s[213] ^ after_pi_s[220];
assign after_theta_s[222] = after_pi_s[222] ^ after_pi_s[225] ^ after_pi_s[232];
assign after_theta_s[234] = after_pi_s[234] ^ after_pi_s[237] ^ after_pi_s[244];
assign after_theta_s[246] = after_pi_s[246] ^ after_pi_s[249] ^ after_pi_s[256];
assign after_theta_s[1] = after_pi_s[1] ^ after_pi_s[4] ^ after_pi_s[11];
assign after_theta_s[13] = after_pi_s[13] ^ after_pi_s[16] ^ after_pi_s[23];
assign after_theta_s[25] = after_pi_s[25] ^ after_pi_s[28] ^ after_pi_s[35];
assign after_theta_s[37] = after_pi_s[37] ^ after_pi_s[40] ^ after_pi_s[47];
assign after_theta_s[49] = after_pi_s[49] ^ after_pi_s[52] ^ after_pi_s[59];
assign after_theta_s[61] = after_pi_s[61] ^ after_pi_s[64] ^ after_pi_s[71];
assign after_theta_s[73] = after_pi_s[73] ^ after_pi_s[76] ^ after_pi_s[83];
assign after_theta_s[85] = after_pi_s[85] ^ after_pi_s[88] ^ after_pi_s[95];
assign after_theta_s[97] = after_pi_s[97] ^ after_pi_s[100] ^ after_pi_s[107];
assign after_theta_s[109] = after_pi_s[109] ^ after_pi_s[112] ^ after_pi_s[119];
assign after_theta_s[121] = after_pi_s[121] ^ after_pi_s[124] ^ after_pi_s[131];
assign after_theta_s[133] = after_pi_s[133] ^ after_pi_s[136] ^ after_pi_s[143];
assign after_theta_s[145] = after_pi_s[145] ^ after_pi_s[148] ^ after_pi_s[155];
assign after_theta_s[157] = after_pi_s[157] ^ after_pi_s[160] ^ after_pi_s[167];
assign after_theta_s[169] = after_pi_s[169] ^ after_pi_s[172] ^ after_pi_s[179];
assign after_theta_s[193] = after_pi_s[193] ^ after_pi_s[196] ^ after_pi_s[203];
assign after_theta_s[205] = after_pi_s[205] ^ after_pi_s[208] ^ after_pi_s[215];
assign after_theta_s[217] = after_pi_s[217] ^ after_pi_s[220] ^ after_pi_s[227];
assign after_theta_s[241] = after_pi_s[241] ^ after_pi_s[244] ^ after_pi_s[251];
assign after_theta_s[253] = after_pi_s[253] ^ after_pi_s[256] ^ after_pi_s[6];
assign after_theta_s[8] = after_pi_s[8] ^ after_pi_s[11] ^ after_pi_s[18];
assign after_theta_s[20] = after_pi_s[20] ^ after_pi_s[23] ^ after_pi_s[30];
assign after_theta_s[32] = after_pi_s[32] ^ after_pi_s[35] ^ after_pi_s[42];
assign after_theta_s[44] = after_pi_s[44] ^ after_pi_s[47] ^ after_pi_s[54];
assign after_theta_s[68] = after_pi_s[68] ^ after_pi_s[71] ^ after_pi_s[78];
assign after_theta_s[80] = after_pi_s[80] ^ after_pi_s[83] ^ after_pi_s[90];
assign after_theta_s[92] = after_pi_s[92] ^ after_pi_s[95] ^ after_pi_s[102];
assign after_theta_s[104] = after_pi_s[104] ^ after_pi_s[107] ^ after_pi_s[114];
assign after_theta_s[116] = after_pi_s[116] ^ after_pi_s[119] ^ after_pi_s[126];
assign after_theta_s[128] = after_pi_s[128] ^ after_pi_s[131] ^ after_pi_s[138];
assign after_theta_s[140] = after_pi_s[140] ^ after_pi_s[143] ^ after_pi_s[150];
assign after_theta_s[164] = after_pi_s[164] ^ after_pi_s[167] ^ after_pi_s[174];
assign after_theta_s[176] = after_pi_s[176] ^ after_pi_s[179] ^ after_pi_s[186];
assign after_theta_s[188] = after_pi_s[188] ^ after_pi_s[191] ^ after_pi_s[198];
assign after_theta_s[200] = after_pi_s[200] ^ after_pi_s[203] ^ after_pi_s[210];
assign after_theta_s[236] = after_pi_s[236] ^ after_pi_s[239] ^ after_pi_s[246];
assign after_theta_s[248] = after_pi_s[248] ^ after_pi_s[251] ^ after_pi_s[1]; 
assign after_theta_s[3] = after_pi_s[3] ^ after_pi_s[6] ^ after_pi_s[13];
assign after_theta_s[15] = after_pi_s[15] ^ after_pi_s[18] ^ after_pi_s[25];
assign after_theta_s[27] = after_pi_s[27] ^ after_pi_s[30] ^ after_pi_s[37];
assign after_theta_s[39] = after_pi_s[39] ^ after_pi_s[42] ^ after_pi_s[49];
assign after_theta_s[63] = after_pi_s[63] ^ after_pi_s[66] ^ after_pi_s[73];
assign after_theta_s[75] = after_pi_s[75] ^ after_pi_s[78] ^ after_pi_s[85];
assign after_theta_s[87] = after_pi_s[87] ^ after_pi_s[90] ^ after_pi_s[97];
assign after_theta_s[99] = after_pi_s[99] ^ after_pi_s[102] ^ after_pi_s[109];
assign after_theta_s[111] = after_pi_s[111] ^ after_pi_s[114] ^ after_pi_s[121];
assign after_theta_s[123] = after_pi_s[123] ^ after_pi_s[126] ^ after_pi_s[133];
assign after_theta_s[135] = after_pi_s[135] ^ after_pi_s[138] ^ after_pi_s[145];
assign after_theta_s[147] = after_pi_s[147] ^ after_pi_s[150] ^ after_pi_s[157];
assign after_theta_s[159] = after_pi_s[159] ^ after_pi_s[162] ^ after_pi_s[169];
assign after_theta_s[171] = after_pi_s[171] ^ after_pi_s[174] ^ after_pi_s[181];
assign after_theta_s[183] = after_pi_s[183] ^ after_pi_s[186] ^ after_pi_s[193];
assign after_theta_s[195] = after_pi_s[195] ^ after_pi_s[198] ^ after_pi_s[205];
assign after_theta_s[207] = after_pi_s[207] ^ after_pi_s[210] ^ after_pi_s[217];
assign after_theta_s[231] = after_pi_s[231] ^ after_pi_s[234] ^ after_pi_s[241];
assign after_theta_s[255] = after_pi_s[255] ^ after_pi_s[1] ^ after_pi_s[8];
assign after_theta_s[10] = after_pi_s[10] ^ after_pi_s[13] ^ after_pi_s[20];
assign after_theta_s[22] = after_pi_s[22] ^ after_pi_s[25] ^ after_pi_s[32];
assign after_theta_s[34] = after_pi_s[34] ^ after_pi_s[37] ^ after_pi_s[44];
assign after_theta_s[46] = after_pi_s[46] ^ after_pi_s[49] ^ after_pi_s[56];
assign after_theta_s[58] = after_pi_s[58] ^ after_pi_s[61] ^ after_pi_s[68];
assign after_theta_s[70] = after_pi_s[70] ^ after_pi_s[73] ^ after_pi_s[80];
assign after_theta_s[82] = after_pi_s[82] ^ after_pi_s[85] ^ after_pi_s[92];
assign after_theta_s[94] = after_pi_s[94] ^ after_pi_s[97] ^ after_pi_s[104];
assign after_theta_s[118] = after_pi_s[118] ^ after_pi_s[121] ^ after_pi_s[128];
assign after_theta_s[142] = after_pi_s[142] ^ after_pi_s[145] ^ after_pi_s[152];
assign after_theta_s[154] = after_pi_s[154] ^ after_pi_s[157] ^ after_pi_s[164];
assign after_theta_s[166] = after_pi_s[166] ^ after_pi_s[169] ^ after_pi_s[176];
assign after_theta_s[178] = after_pi_s[178] ^ after_pi_s[181] ^ after_pi_s[188];
assign after_theta_s[190] = after_pi_s[190] ^ after_pi_s[193] ^ after_pi_s[200];
assign after_theta_s[202] = after_pi_s[202] ^ after_pi_s[205] ^ after_pi_s[212];
assign after_theta_s[214] = after_pi_s[214] ^ after_pi_s[217] ^ after_pi_s[224];
assign after_theta_s[226] = after_pi_s[226] ^ after_pi_s[229] ^ after_pi_s[236];
assign after_theta_s[250] = after_pi_s[250] ^ after_pi_s[253] ^ after_pi_s[3];
assign after_theta_s[5] = after_pi_s[5] ^ after_pi_s[8] ^ after_pi_s[15];
assign after_theta_s[17] = after_pi_s[17] ^ after_pi_s[20] ^ after_pi_s[27];
assign after_theta_s[29] = after_pi_s[29] ^ after_pi_s[32] ^ after_pi_s[39];
assign after_theta_s[41] = after_pi_s[41] ^ after_pi_s[44] ^ after_pi_s[51];
assign after_theta_s[53] = after_pi_s[53] ^ after_pi_s[56] ^ after_pi_s[63];
assign after_theta_s[77] = after_pi_s[77] ^ after_pi_s[80] ^ after_pi_s[87];
assign after_theta_s[89] = after_pi_s[89] ^ after_pi_s[92] ^ after_pi_s[99];
assign after_theta_s[101] = after_pi_s[101] ^ after_pi_s[104] ^ after_pi_s[111];
assign after_theta_s[113] = after_pi_s[113] ^ after_pi_s[116] ^ after_pi_s[123];
assign after_theta_s[125] = after_pi_s[125] ^ after_pi_s[128] ^ after_pi_s[135];
assign after_theta_s[137] = after_pi_s[137] ^ after_pi_s[140] ^ after_pi_s[147];
assign after_theta_s[149] = after_pi_s[149] ^ after_pi_s[152] ^ after_pi_s[159];
assign after_theta_s[173] = after_pi_s[173] ^ after_pi_s[176] ^ after_pi_s[183];
assign after_theta_s[185] = after_pi_s[185] ^ after_pi_s[188] ^ after_pi_s[195];
assign after_theta_s[197] = after_pi_s[197] ^ after_pi_s[200] ^ after_pi_s[207];
assign after_theta_s[209] = after_pi_s[209] ^ after_pi_s[212] ^ after_pi_s[219];
assign after_theta_s[221] = after_pi_s[221] ^ after_pi_s[224] ^ after_pi_s[231];
assign after_theta_s[233] = after_pi_s[233] ^ after_pi_s[236] ^ after_pi_s[243];


// Chi step
assign round_o[254:0] = after_theta_s[254:0] ^   ((~after_theta_s[255:1]) & after_theta_s[256:2]);
assign round_o[255]   = after_theta_s[255]   ^   ((~after_theta_s[256])   & after_theta_s[0]);
assign round_o[256]   = after_theta_s[256]   ^   ((~after_theta_s[0])     & after_theta_s[1]);


endmodule



